library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity ram_2k is
    Port (
       clk   : in  std_logic;
       rst   : in  std_logic;
       cs    : in  std_logic;
       rw    : in  std_logic;
       addr  : in  std_logic_vector (10 downto 0);
       rdata : out std_logic_vector (7 downto 0);
       wdata : in  std_logic_vector (7 downto 0)
    );
end ram_2k;

architecture rtl of ram_2k is


signal we : std_logic;
signal dp : std_logic;

begin

  ROM : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do     => rdata,
	  dop(0) => dp,
	  addr   => addr,
	  clk    => clk,
	  di     => wdata,
	  dip(0) => dp,
	  en     => cs,
	  ssr    => rst,
	  we     => we
	);

my_ram_2k : process ( rw )
begin
	 we    <= not rw;
end process;

end architecture rtl;

